package test_pkg;

  import i2c_pkg::*;

  include "base_test.sv";
  include "i2c_standard_test.sv";
  include "i2c_fast_test.sv";
  include "i2c_fast_plus_test.sv";

endpackage