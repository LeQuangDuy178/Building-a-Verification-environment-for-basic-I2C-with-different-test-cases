package i2c_pkg;

    `include "packet.sv"
    `include "stimulus.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "environment.sv"

endpackage